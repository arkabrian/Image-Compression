library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity downscale_tb is
end entity downscale_tb;

architecture rtl of downscale_tb is

begin

  

end architecture;